`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/25/2016 12:41:21 PM
// Design Name: 
// Module Name: Checking_nbits
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// Check if one-bit input is correct
module Checking_1bit(
    output correct,
    output checking_done,
    output [1:0] led_pressed,
    input clock,
    input right_pressed,
    input left_pressed,
    input bit_gen      // bit generated by random number generator
    );

reg correct_reg;
reg [1:0] led_pressed_reg;
reg input_bit;
reg done;

assign correct = correct_reg;
assign led_pressed = led_pressed_reg;
assign checking_done = done;

always @(posedge clock)
    begin
    if(right_pressed==1) begin
        input_bit <= 1;
        led_pressed_reg = 2'b01;
        done = 0;
        end        
    else if(left_pressed==1) begin
        input_bit = 0;
        led_pressed_reg = 2'b10;
        done = 0;
        end
    else begin
        led_pressed_reg = 2'b00;
        done = 0;
        end
        
    if(input_bit==bit_gen)  begin
        correct_reg <= 1;
        done <= 1;
        end
    else begin
        correct_reg <= 0;
        done <= 1;
        end
    end   

endmodule

//--------------------------------------------------------------
// Check if n-bit input sequence is correct
module Checking_nbits(      
    output correct,
    output checking_done,
    output [1:0] led_pressed_n,
    output [3:0] index,
    input clock,
    input right_pressed,
    input left_pressed,
    input enable,
    input [2:0] bit_count,  // number of bits in sequence  
    input [7:0] bit_gen_sequence   // bit sequence generated by random number generator
    );
    
reg correct_stat;    
reg correct_reg;
reg [1:0] led_reg;
reg done;
wire temp;
wire checking_done_temp;
wire [1:0] led_pressed;
reg checking_temp_reg;
reg [3:0] i;
reg state;

assign correct = correct_reg;
assign checking_done = done;
assign led_pressed_n = led_reg;
assign index = i;

initial begin   
    i<= 0;
    correct_stat <= 1;
    correct_reg <= 0;
    done <= 0;
    checking_temp_reg <= 0;
    state <= 0;
    end
    
Checking_1bit Check(temp, checking_done_temp, led_pressed, clock, right_pressed, left_pressed, bit_gen_sequence[i]);

always @(posedge clock) begin
    led_reg = led_pressed;
    if(enable == 1) begin
    if(done == 1)   i = i;
    else begin
        case(state)
            0: begin
                if(right_pressed || left_pressed) begin
                    checking_temp_reg = checking_done_temp;
                    if(checking_temp_reg == 1)  begin
                        correct_stat = temp;
                        state <= 1;
                        end
                    else state <= 0;
                    end
                else state <= 0;
                end
            1: begin
                if((correct_stat == 0)|| (i>=bit_count)) begin
                    correct_reg = correct_stat;
                    done = 1;
                    i = i;
                    end
                else if((correct_stat == 1)&&(i<bit_count)) begin
                    done = 0;
                    i = i + 1;
                    state <= 0;
                    end
                end
            endcase
        end
        end
    else begin
        i<= 0;
        correct_stat <= 1;
        correct_reg <= 0;
        done <= 0;
        checking_temp_reg <= 0;
        state <= 0;
        end
    end
        
                
    
endmodule
