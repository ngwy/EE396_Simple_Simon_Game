`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/25/2016 12:41:21 PM
// Design Name: 
// Module Name: Checking_nbits
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// Check if one-bit input is correct
module Checking_1bit(
    output          correct,
    output [1:0]    led_pressed,
    input           clock,
    input           right_pressed,
    input           left_pressed,
    input           enable,
    input           bit_gen      // bit generated by random number generator
    );

reg         correct_reg;
reg  [1:0]  led_pressed_reg;

assign      correct         = correct_reg;
assign      led_pressed     = led_pressed_reg;

always @(posedge clock) begin
    if (enable) begin
        if (right_pressed == 1) begin
            led_pressed_reg     <= 0'b01;
            if (bit_gen == 1)   correct_reg <= 1;
            else                correct_reg <= 0;
            end
        else if (left_pressed == 1) begin
            led_pressed_reg     <= 0'b10;
            if (bit_gen == 0)   correct_reg <= 1;
            else                correct_reg <= 0;
            end
        else    led_pressed_reg <= 0'b00;
        end
    else
        led_pressed_reg         <= 0'b00;
    end

endmodule

//--------------------------------------------------------------
// Check if n-bit input sequence is correct
//module Checking_nbits(      
//    output          correct,
//    output          checking_done,
//    output [1:0]    led_pressed_n,
//    output [3:0]    index,
//    input           clock,
//    input           right_pressed,
//    input           left_pressed,
//    input           enable,
//    input  [2:0]    bit_count,  // number of bits in sequence  
//    input  [7:0]    bit_gen_sequence   // bit sequence generated by random number generator
//    );

//wire        temp;
//wire        checking_done_temp;
//wire [1:0]  led_pressed;

//reg  [1:0]  led_reg; 
//reg  [3:0]  i;   
//reg         bit_enable;
//reg         checking_temp_reg;
//reg         correct_stat;    
//reg         correct_reg;
//reg         done;
//reg         state;

//assign      correct         = correct_reg;
//assign      checking_done   = done;
//assign      led_pressed_n   = led_reg;
//assign      index           = i;

//initial begin   
//    i                   <= 0;
//    bit_enable          <= 0;
//    correct_stat        <= 0;
//    correct_reg         <= 0;
//    done                <= 0;
//    end

//Checking_1bit   Check(temp, led_pressed, clock, right_pressed, left_pressed, bit_enable, bit_gen_sequence[i]);

//always @(posedge clock) begin
//    led_reg <= led_pressed;
//    if  (enable == 1) begin
//        if (i <= bit_count) begin
//            bit_enable <= 1;
//            if (right_pressed == 1 || left_pressed == 1) begin
//                correct_stat    <= temp;
//                if (correct_stat == 0) begin
//                    correct_reg <= 0;
//                    bit_enable  <= 0;
//                    done = 1;
//                    end
//                else begin
//                    done <= 0;
//                    i <= i + 1;
//                    end
//                end
//            else   begin
//                done <= 0;
//                i <= i;
//                end
//            end
//        else begin
//            correct_reg = 1;
//            bit_enable  = 0;
//            done        = 1;
//            end      
                    
            
//        end
//    else begin
//     i                   = 0;
//    bit_enable          = 0;
//    correct_stat        = 0;
//    correct_reg         = 0;
//    done                = 0;
            
//    end
//     end   
                
//endmodule
